`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/28/2023 01:32:58 PM
// Design Name: 
// Module Name: register
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module RF(A, B, SA, SB, D, DA, W, rst, clk);
output [3:0]A; // A bus
output [3:0]B; // B bus
input SA; // Select A - A Address
input SB; // Select B - B Address
input [3:0]D; // Data input
input DA; // Data destination address
input W; // write enable
input rst; // positive logic asynchronous reset
input clk;
wire [1:0]load_enable;
wire [3:0]R00, R01;

Decoder1to2 decoder (load_enable, DA, W);
RegisterNbit reg00 (D,R00,load_enable[0], rst, clk); //D-in, R00-out
RegisterNbit reg01 (D,R01,load_enable[1], rst, clk);
Mux2to1Nbit muxA (A,R00, R01, SA);
Mux2to1Nbit muxB (B,R00, R01,SB);
endmodule

module RegisterNbit(D, Q, L, R, clock);
parameter N = 4; // number of bits
output reg [N-1:0]Q; // registered output
input [N-1:0]D; // data input
input L; // load enable
input R; // positive logic asynchronous reset
input clock; // positive edge clock

always @(posedge clock or posedge R) begin
if(R)
Q<=0;
else if(L)
Q<=D;
else
Q<=Q;

end
endmodule

module Decoder1to2(m, S, en);
input S; // select
input en; // enable (positive logic)
output [1:0]m; // 32 minterms
assign m[0] = ~S&en;
assign m[1] = S&en;
endmodule

module Mux2to1Nbit(o, i1,i2, s);
input [3:0] i1,i2;
input s;
output reg [3:0] o;
always @(s or i1 or i2)
begin
case (s)
1'b0 : o = i1;
1'b1 : o = i2;
default : o = 4'b0;
endcase
end
endmodule
